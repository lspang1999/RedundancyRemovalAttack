
module c880
(
  N1,
  N8,
  N13,
  N17,
  N26,
  N29,
  N36,
  N42,
  N51,
  N55,
  N59,
  N68,
  N72,
  N73,
  N74,
  N75,
  N80,
  N85,
  N86,
  N87,
  N88,
  N89,
  N90,
  N91,
  N96,
  N101,
  N106,
  N111,
  N116,
  N121,
  N126,
  N130,
  N135,
  N138,
  N143,
  N146,
  N149,
  N152,
  N153,
  N156,
  N159,
  N165,
  N171,
  N177,
  N183,
  N189,
  N195,
  N201,
  N207,
  N210,
  N219,
  N228,
  N237,
  N246,
  N255,
  N259,
  N260,
  N261,
  N267,
  N268,
  N388,
  N389,
  N390,
  N391,
  N418,
  N419,
  N420,
  N421,
  N422,
  N423,
  N446,
  N447,
  N448,
  N449,
  N450,
  N767,
  N768,
  N850,
  N863,
  N864,
  N865,
  N866,
  N874,
  N878,
  N879,
  N880,
  keyInput0,
  keyInput1,
  keyInput2,
  keyInput3,
  keyInput4,
  keyInput5,
  keyInput6,
  keyInput7,
  keyInput8,
  keyInput9,
  keyInput10,
  keyInput11,
  keyInput12,
  keyInput13,
  keyInput14,
  keyInput15,
  keyInput16,
  keyInput17,
  keyInput18
);

  input N1;input N8;input N13;input N17;input N26;input N29;input N36;input N42;input N51;input N55;input N59;input N68;input N72;input N73;input N74;input N75;input N80;input N85;input N86;input N87;input N88;input N89;input N90;input N91;input N96;input N101;input N106;input N111;input N116;input N121;input N126;input N130;input N135;input N138;input N143;input N146;input N149;input N152;input N153;input N156;input N159;input N165;input N171;input N177;input N183;input N189;input N195;input N201;input N207;input N210;input N219;input N228;input N237;input N246;input N255;input N259;input N260;input N261;input N267;input N268;output N388;output N389;output N390;output N391;output N418;output N419;output N420;output N421;output N422;output N423;output N446;output N447;output N448;output N449;output N450;output N767;output N768;output N850;output N863;output N864;output N865;output N866;output N874;output N878;output N879;output N880;wire N269;wire N270;wire N273;wire N276;wire N279;wire N280;wire N284;wire N285;wire N286;wire N287;wire N290;wire N291;wire N292;wire N293;wire N294;wire N295;wire N296;wire N297;wire N298;wire N301;wire N302;wire N303;wire N304;wire N305;wire N306;wire N307;wire N308;wire N309;wire N310;wire N316;wire N317;wire N318;wire N319;wire N322;wire N323;wire N324;wire N325;wire N326;wire N327;wire N328;wire N329;wire N330;wire N331;wire N332;wire N333;wire N334;wire N335;wire N336;wire N337;wire N338;wire N339;wire N340;wire N341;wire N342;wire N343;wire N344;wire N345;wire N346;wire N347;wire N348;wire N349;wire N350;wire N351;wire N352;wire N353;wire N354;wire N355;wire N356;wire N357;wire N360;wire N363;wire N366;wire N369;wire N375;wire N376;wire N379;wire N382;wire N385;wire N392;wire N393;wire N399;wire N400;wire N401;wire N402;wire N403;wire N404;wire N405;wire N406;wire N407;wire N408;wire N409;wire N410;wire N411;wire N412;wire N413;wire N414;wire N415;wire N416;wire N417;wire N424;wire N425;wire N426;wire N427;wire N432;wire N437;wire N442;wire N443;wire N444;wire N445;wire N451;wire N460;wire N463;wire N466;wire N475;wire N476;wire N477;wire N478;wire N479;wire N480;wire N481;wire N482;wire N483;wire N488;wire N489;wire N490;wire N491;wire N492;wire N495;wire N498;wire N499;wire N500;wire N501;wire N502;wire N503;wire N504;wire N505;wire N506;wire N507;wire N508;wire N509;wire N510;wire N511;wire N512;wire N513;wire N514;wire N515;wire N516;wire N517;wire N518;wire N519;wire N520;wire N521;wire N522;wire N523;wire N524;wire N525;wire N526;wire N527;wire N528;wire N529;wire N530;wire N533;wire N536;wire N537;wire N538;wire N539;wire N540;wire N541;wire N542;wire N543;wire N544;wire N547;wire N550;wire N551;wire N552;wire N553;wire N557;wire N561;wire N565;wire N569;wire N573;wire N577;wire N581;wire N585;wire N586;wire N587;wire N588;wire N589;wire N590;wire N593;wire N596;wire N597;wire N600;wire N605;wire N606;wire N609;wire N615;wire N616;wire N619;wire N624;wire N625;wire N628;wire N631;wire N632;wire N635;wire N640;wire N641;wire N644;wire N650;wire N651;wire N654;wire N659;wire N660;wire N661;wire N662;wire N665;wire N669;wire N670;wire N673;wire N677;wire N678;wire N682;wire N686;wire N687;wire N692;wire N696;wire N697;wire N700;wire N704;wire N705;wire N708;wire N712;wire N713;wire N717;wire N721;wire N722;wire N727;wire N731;wire N732;wire N733;wire N734;wire N735;wire N736;wire N737;wire N738;wire N739;wire N740;wire N741;wire N742;wire N743;wire N744;wire N745;wire N746;wire N747;wire N748;wire N749;wire N750;wire N751;wire N752;wire N753;wire N754;wire N755;wire N756;wire N757;wire N758;wire N759;wire N760;wire N761;wire N762;wire N763;wire N764;wire N765;wire N766;wire N769;wire N770;wire N771;wire N772;wire N773;wire N777;wire N778;wire N781;wire N782;wire N785;wire N786;wire N787;wire N788;wire N789;wire N790;wire N791;wire N792;wire N793;wire N794;wire N795;wire N796;wire N802;wire N803;wire N804;wire N805;wire N806;wire N807;wire N808;wire N809;wire N810;wire N811;wire N812;wire N813;wire N814;wire N815;wire N819;wire N822;wire N825;wire N826;wire N827;wire N828;wire N829;wire N830;wire N831;wire N832;wire N833;wire N834;wire N835;wire N836;wire N837;wire N838;wire N839;wire N840;wire N841;wire N842;wire N843;wire N844;wire N845;wire N846;wire N847;wire N848;wire N849;wire N851;wire N852;wire N853;wire N854;wire N855;wire N856;wire N857;wire N858;wire N859;wire N860;wire N861;wire N862;wire N867;wire N868;wire N869;wire N870;wire N871;wire N872;wire N873;wire N875;wire N876;wire N877;wire keyWire0;input keyInput0;wire keyWire1;input keyInput1;wire keyWire2;input keyInput2;wire keyWire3;input keyInput3;wire keyWire4;input keyInput4;wire keyWire5;input keyInput5;wire keyWire6;input keyInput6;wire keyWire7;input keyInput7;wire keyWire8;input keyInput8;wire keyWire9;input keyInput9;wire keyWire10;input keyInput10;wire keyWire11;input keyInput11;wire keyWire12;input keyInput12;wire keyWire13;input keyInput13;wire keyWire14;input keyInput14;wire keyWire15;input keyInput15;wire keyWire16;input keyInput16;wire keyWire17;input keyInput17;wire keyWire18;input keyInput18;

  nand
  NAND4_1
  (
    N269,
    N1,
    N8,
    N13,
    N17
  );


  nand
  NAND4_2
  (
    N270,
    N1,
    N26,
    N13,
    N17
  );


  and
  AND3_3
  (
    N273,
    N29,
    N36,
    N42
  );


  and
  AND3_4
  (
    N276,
    N1,
    N26,
    N51
  );


  nand
  NAND4_6
  (
    N280,
    N1,
    N8,
    N13,
    N55
  );


  nand
  NAND4_7
  (
    N284,
    N59,
    N42,
    N68,
    N72
  );


  nand
  NAND2_8
  (
    N285,
    N29,
    N68
  );


  nand
  NAND3_9
  (
    N286,
    N59,
    N68,
    N74
  );


  and
  AND3_10
  (
    N287,
    N29,
    N75,
    N80
  );


  and
  AND3_11
  (
    N290,
    N29,
    N75,
    N42
  );


  and
  AND3_12
  (
    N291,
    N29,
    N36,
    N80
  );


  and
  AND3_13
  (
    N292,
    N29,
    N36,
    N42
  );


  and
  AND3_14
  (
    N293,
    N59,
    N75,
    N80
  );


  and
  AND3_15
  (
    N294,
    N59,
    N75,
    N42
  );


  and
  AND3_16
  (
    N295,
    N59,
    N36,
    N80
  );


  and
  AND3_17
  (
    N296,
    N59,
    N36,
    N42
  );


  and
  AND2_18
  (
    N297,
    N85,
    N86
  );


  or
  OR2_19
  (
    N298,
    N87,
    N88
  );


  nand
  NAND2_20
  (
    N301,
    N91,
    N96
  );


  or
  OR2_21
  (
    N302,
    N91,
    N96
  );


  or
  OR2_23
  (
    N304,
    N101,
    N106
  );


  or
  OR2_25
  (
    N306,
    N111,
    N116
  );


  nand
  NAND2_26
  (
    N307,
    N121,
    N126
  );


  or
  OR2_27
  (
    N308,
    N121,
    N126
  );


  and
  AND2_28
  (
    N309,
    N8,
    N138
  );


  not
  NOT1_29
  (
    N310,
    N268
  );


  and
  AND2_30
  (
    N316,
    N51,
    N138
  );


  and
  AND2_31
  (
    N317,
    N17,
    N138
  );


  and
  AND2_32
  (
    N318,
    N152,
    N138
  );


  nand
  NAND2_33
  (
    N319,
    N59,
    N156
  );


  nor
  NOR2_34
  (
    N322,
    N17,
    N42
  );


  and
  AND2_35
  (
    N323,
    N17,
    N42
  );


  nand
  NAND2_36
  (
    N324,
    N159,
    N165
  );


  or
  OR2_37
  (
    N325,
    N159,
    N165
  );


  nand
  NAND2_38
  (
    N326,
    N171,
    N177
  );


  or
  OR2_39
  (
    N327,
    N171,
    N177
  );


  nand
  NAND2_40
  (
    N328,
    N183,
    N189
  );


  or
  OR2_41
  (
    N329,
    N183,
    N189
  );


  nand
  NAND2_42
  (
    N330,
    N195,
    N201
  );


  or
  OR2_43
  (
    N331,
    N195,
    N201
  );


  and
  AND2_44
  (
    N332,
    N210,
    N91
  );


  and
  AND2_45
  (
    N333,
    N210,
    N96
  );


  and
  AND2_46
  (
    N334,
    N210,
    N101
  );


  and
  AND2_47
  (
    N335,
    N210,
    N106
  );


  and
  AND2_48
  (
    N336,
    N210,
    N111
  );


  and
  AND2_49
  (
    N337,
    N255,
    N259
  );


  and
  AND2_50
  (
    N338,
    N210,
    N116
  );


  and
  AND2_51
  (
    N339,
    N255,
    N260
  );


  and
  AND2_52
  (
    N340,
    N210,
    N121
  );


  and
  AND2_53
  (
    N341,
    N255,
    N267
  );


  not
  NOT1_54
  (
    N342,
    N269
  );


  not
  NOT1_55
  (
    N343,
    N273
  );


  or
  OR2_56
  (
    N344,
    N270,
    N273
  );


  not
  NOT1_57
  (
    N345,
    N276
  );


  not
  NOT1_58
  (
    N346,
    N276
  );


  not
  NOT1_59
  (
    N347,
    N279
  );


  nor
  NOR2_60
  (
    N348,
    N280,
    N284
  );


  or
  OR2_61
  (
    N349,
    N280,
    N285
  );


  or
  OR2_62
  (
    N350,
    N280,
    N286
  );


  not
  NOT1_63
  (
    N351,
    N293
  );


  not
  NOT1_64
  (
    N352,
    N294
  );


  not
  NOT1_65
  (
    N353,
    N295
  );


  not
  NOT1_66
  (
    N354,
    N296
  );


  and
  AND2_68
  (
    N356,
    N90,
    N298
  );


  nand
  NAND2_69
  (
    N357,
    N301,
    N302
  );


  nand
  NAND2_70
  (
    N360,
    N303,
    N304
  );


  nand
  NAND2_71
  (
    N363,
    N305,
    N306
  );


  nand
  NAND2_72
  (
    N366,
    N307,
    N308
  );


  not
  NOT1_73
  (
    N369,
    N310
  );


  nor
  NOR2_74
  (
    N375,
    N322,
    N323
  );


  nand
  NAND2_75
  (
    N376,
    N324,
    N325
  );


  nand
  NAND2_76
  (
    N379,
    N326,
    N327
  );


  nand
  NAND2_77
  (
    N382,
    N328,
    N329
  );


  nand
  NAND2_78
  (
    N385,
    N330,
    N331
  );


  buf
  BUFF1_79
  (
    N388,
    N290
  );


  buf
  BUFF1_81
  (
    N390,
    N292
  );


  buf
  BUFF1_82
  (
    N391,
    N297
  );


  or
  OR2_83
  (
    N392,
    N270,
    N343
  );


  not
  NOT1_84
  (
    N393,
    N345
  );


  not
  NOT1_85
  (
    N399,
    N346
  );


  and
  AND2_86
  (
    N400,
    N348,
    N73
  );


  not
  NOT1_87
  (
    N401,
    N349
  );


  not
  NOT1_88
  (
    N402,
    N350
  );


  not
  NOT1_89
  (
    N403,
    N355
  );


  not
  NOT1_90
  (
    N404,
    N357
  );


  not
  NOT1_91
  (
    N405,
    N360
  );


  and
  AND2_92
  (
    N406,
    N357,
    N360
  );


  not
  NOT1_93
  (
    N407,
    N363
  );


  not
  NOT1_94
  (
    N408,
    N366
  );


  and
  AND2_95
  (
    N409,
    N363,
    N366
  );


  nand
  NAND2_96
  (
    N410,
    N347,
    N352
  );


  not
  NOT1_97
  (
    N411,
    N376
  );


  not
  NOT1_98
  (
    N412,
    N379
  );


  and
  AND2_99
  (
    N413,
    N376,
    N379
  );


  not
  NOT1_100
  (
    N414,
    N382
  );


  not
  NOT1_101
  (
    N415,
    N385
  );


  and
  AND2_102
  (
    N416,
    N382,
    N385
  );


  and
  AND2_103
  (
    N417,
    N210,
    N369
  );


  buf
  BUFF1_104
  (
    N418,
    N342
  );


  buf
  BUFF1_105
  (
    N419,
    N344
  );


  buf
  BUFF1_106
  (
    N420,
    N351
  );


  buf
  BUFF1_107
  (
    N421,
    N353
  );


  buf
  BUFF1_108
  (
    N422,
    N354
  );


  not
  NOT1_110
  (
    N424,
    N400
  );


  and
  AND2_111
  (
    N425,
    N404,
    N405
  );


  and
  AND2_112
  (
    N426,
    N407,
    N408
  );


  and
  AND3_113
  (
    N427,
    N319,
    N393,
    N55
  );


  and
  AND3_114
  (
    N432,
    N393,
    N17,
    N287
  );


  nand
  NAND3_115
  (
    N437,
    N393,
    N287,
    N55
  );


  nand
  NAND4_116
  (
    N442,
    N375,
    N59,
    N156,
    N393
  );


  nand
  NAND3_117
  (
    N443,
    N393,
    N319,
    N17
  );


  and
  AND2_118
  (
    N444,
    N411,
    N412
  );


  and
  AND2_119
  (
    N445,
    N414,
    N415
  );


  buf
  BUFF1_120
  (
    N446,
    N392
  );


  buf
  BUFF1_121
  (
    N447,
    N399
  );


  buf
  BUFF1_122
  (
    N448,
    N401
  );


  buf
  BUFF1_123
  (
    N449,
    N402
  );


  buf
  BUFF1_124
  (
    N450,
    N403
  );


  not
  NOT1_125
  (
    N451,
    N424
  );


  nor
  NOR2_126
  (
    N460,
    N406,
    N425
  );


  nor
  NOR2_127
  (
    N463,
    N409,
    N426
  );


  nand
  NAND2_128
  (
    N466,
    N442,
    N410
  );


  and
  AND2_129
  (
    N475,
    N143,
    N427
  );


  and
  AND2_130
  (
    N476,
    N310,
    N432
  );


  and
  AND2_131
  (
    N477,
    N146,
    N427
  );


  and
  AND2_132
  (
    N478,
    N310,
    N432
  );


  and
  AND2_133
  (
    N479,
    N149,
    N427
  );


  and
  AND2_134
  (
    N480,
    N310,
    N432
  );


  and
  AND2_135
  (
    N481,
    N153,
    N427
  );


  and
  AND2_136
  (
    N482,
    N310,
    N432
  );


  nand
  NAND2_137
  (
    N483,
    N443,
    N1
  );


  or
  OR2_138
  (
    N488,
    N369,
    N437
  );


  or
  OR2_139
  (
    N489,
    N369,
    N437
  );


  or
  OR2_140
  (
    N490,
    N369,
    N437
  );


  or
  OR2_141
  (
    N491,
    N369,
    N437
  );


  nor
  NOR2_142
  (
    N492,
    N413,
    N444
  );


  nor
  NOR2_143
  (
    N495,
    N416,
    N445
  );


  nand
  NAND2_144
  (
    N498,
    N130,
    N460
  );


  or
  OR2_145
  (
    N499,
    N130,
    N460
  );


  nand
  NAND2_146
  (
    N500,
    N463,
    N135
  );


  or
  OR2_147
  (
    N501,
    N463,
    N135
  );


  and
  AND2_148
  (
    N502,
    N91,
    N466
  );


  nor
  NOR2_149
  (
    N503,
    N475,
    N476
  );


  and
  AND2_150
  (
    N504,
    N96,
    N466
  );


  nor
  NOR2_151
  (
    N505,
    N477,
    N478
  );


  and
  AND2_152
  (
    N506,
    N101,
    N466
  );


  nor
  NOR2_153
  (
    N507,
    N479,
    N480
  );


  and
  AND2_154
  (
    N508,
    N106,
    N466
  );


  nor
  NOR2_155
  (
    N509,
    N481,
    N482
  );


  and
  AND2_156
  (
    N510,
    N143,
    N483
  );


  and
  AND2_158
  (
    N512,
    N146,
    N483
  );


  and
  AND2_159
  (
    N513,
    N116,
    N466
  );


  and
  AND2_160
  (
    N514,
    N149,
    N483
  );


  and
  AND2_161
  (
    N515,
    N121,
    N466
  );


  and
  AND2_162
  (
    N516,
    N153,
    N483
  );


  nand
  NAND2_164
  (
    N518,
    N130,
    N492
  );


  or
  OR2_165
  (
    N519,
    N130,
    N492
  );


  nand
  NAND2_166
  (
    N520,
    N495,
    N207
  );


  or
  OR2_167
  (
    N521,
    N495,
    N207
  );


  and
  AND2_168
  (
    N522,
    N451,
    N159
  );


  and
  AND2_169
  (
    N523,
    N451,
    N165
  );


  and
  AND2_171
  (
    N525,
    N451,
    N177
  );


  and
  AND2_172
  (
    N526,
    N451,
    N183
  );


  nand
  NAND2_173
  (
    N527,
    N451,
    N189
  );


  nand
  NAND2_174
  (
    N528,
    N451,
    N195
  );


  nand
  NAND2_175
  (
    N529,
    N451,
    N201
  );


  nand
  NAND2_176
  (
    N530,
    N498,
    N499
  );


  nand
  NAND2_177
  (
    N533,
    N500,
    N501
  );


  nor
  NOR2_178
  (
    N536,
    N309,
    N502
  );


  nor
  NOR2_179
  (
    N537,
    N316,
    N504
  );


  nor
  NOR2_180
  (
    N538,
    N317,
    N506
  );


  nor
  NOR2_182
  (
    N540,
    N510,
    N511
  );


  nor
  NOR2_183
  (
    N541,
    N512,
    N513
  );


  nor
  NOR2_184
  (
    N542,
    N514,
    N515
  );


  nor
  NOR2_185
  (
    N543,
    N516,
    N517
  );


  nand
  NAND2_186
  (
    N544,
    N518,
    N519
  );


  nand
  NAND2_187
  (
    N547,
    N520,
    N521
  );


  not
  NOT1_188
  (
    N550,
    N530
  );


  not
  NOT1_189
  (
    N551,
    N533
  );


  and
  AND2_190
  (
    N552,
    N530,
    N533
  );


  nand
  NAND2_191
  (
    N553,
    N536,
    N503
  );


  nand
  NAND2_192
  (
    N557,
    N537,
    N505
  );


  nand
  NAND2_193
  (
    N561,
    N538,
    N507
  );


  nand
  NAND2_194
  (
    N565,
    N539,
    N509
  );


  nand
  NAND2_195
  (
    N569,
    N488,
    N540
  );


  nand
  NAND2_196
  (
    N573,
    N489,
    N541
  );


  nand
  NAND2_197
  (
    N577,
    N490,
    N542
  );


  nand
  NAND2_198
  (
    N581,
    N491,
    N543
  );


  not
  NOT1_199
  (
    N585,
    N544
  );


  not
  NOT1_200
  (
    N586,
    N547
  );


  and
  AND2_201
  (
    N587,
    N544,
    N547
  );


  and
  AND2_202
  (
    N588,
    N550,
    N551
  );


  and
  AND2_203
  (
    N589,
    N585,
    N586
  );


  or
  OR2_205
  (
    N593,
    N553,
    N159
  );


  and
  AND2_206
  (
    N596,
    N246,
    N553
  );


  nand
  NAND2_207
  (
    N597,
    N557,
    N165
  );


  or
  OR2_208
  (
    N600,
    N557,
    N165
  );


  and
  AND2_209
  (
    N605,
    N246,
    N557
  );


  nand
  NAND2_210
  (
    N606,
    N561,
    N171
  );


  or
  OR2_211
  (
    N609,
    N561,
    N171
  );


  and
  AND2_212
  (
    N615,
    N246,
    N561
  );


  nand
  NAND2_213
  (
    N616,
    N565,
    N177
  );


  or
  OR2_214
  (
    N619,
    N565,
    N177
  );


  and
  AND2_215
  (
    N624,
    N246,
    N565
  );


  nand
  NAND2_216
  (
    N625,
    N569,
    N183
  );


  or
  OR2_217
  (
    N628,
    N569,
    N183
  );


  and
  AND2_218
  (
    N631,
    N246,
    N569
  );


  nand
  NAND2_219
  (
    N632,
    N573,
    N189
  );


  or
  OR2_220
  (
    N635,
    N573,
    N189
  );


  and
  AND2_221
  (
    N640,
    N246,
    N573
  );


  nand
  NAND2_222
  (
    N641,
    N577,
    N195
  );


  and
  AND2_224
  (
    N650,
    N246,
    N577
  );


  nand
  NAND2_225
  (
    N651,
    N581,
    N201
  );


  or
  OR2_226
  (
    N654,
    N581,
    N201
  );


  nor
  NOR2_228
  (
    N660,
    N552,
    N588
  );


  nor
  NOR2_229
  (
    N661,
    N587,
    N589
  );


  not
  NOT1_230
  (
    N662,
    N590
  );


  and
  AND2_231
  (
    N665,
    N593,
    N590
  );


  nor
  NOR2_232
  (
    N669,
    N596,
    N522
  );


  not
  NOT1_233
  (
    N670,
    N597
  );


  and
  AND2_234
  (
    N673,
    N600,
    N597
  );


  nor
  NOR2_235
  (
    N677,
    N605,
    N523
  );


  not
  NOT1_236
  (
    N678,
    N606
  );


  and
  AND2_237
  (
    N682,
    N609,
    N606
  );


  nor
  NOR2_238
  (
    N686,
    N615,
    N524
  );


  not
  NOT1_239
  (
    N687,
    N616
  );


  and
  AND2_240
  (
    N692,
    N619,
    N616
  );


  nor
  NOR2_241
  (
    N696,
    N624,
    N525
  );


  not
  NOT1_242
  (
    N697,
    N625
  );


  and
  AND2_243
  (
    N700,
    N628,
    N625
  );


  nor
  NOR2_244
  (
    N704,
    N631,
    N526
  );


  not
  NOT1_245
  (
    N705,
    N632
  );


  and
  AND2_246
  (
    N708,
    N635,
    N632
  );


  nor
  NOR2_247
  (
    N712,
    N337,
    N640
  );


  not
  NOT1_248
  (
    N713,
    N641
  );


  nor
  NOR2_250
  (
    N721,
    N339,
    N650
  );


  not
  NOT1_251
  (
    N722,
    N651
  );


  and
  AND2_252
  (
    N727,
    N654,
    N651
  );


  nor
  NOR2_253
  (
    N731,
    N341,
    N659
  );


  nand
  NAND2_254
  (
    N732,
    N654,
    N261
  );


  nand
  NAND3_255
  (
    N733,
    N644,
    N654,
    N261
  );


  nand
  NAND4_256
  (
    N734,
    N635,
    N644,
    N654,
    N261
  );


  not
  NOT1_257
  (
    N735,
    N662
  );


  and
  AND2_258
  (
    N736,
    N228,
    N665
  );


  and
  AND2_259
  (
    N737,
    N237,
    N662
  );


  not
  NOT1_260
  (
    N738,
    N670
  );


  and
  AND2_261
  (
    N739,
    N228,
    N673
  );


  and
  AND2_262
  (
    N740,
    N237,
    N670
  );


  not
  NOT1_263
  (
    N741,
    N678
  );


  and
  AND2_264
  (
    N742,
    N228,
    N682
  );


  and
  AND2_265
  (
    N743,
    N237,
    N678
  );


  not
  NOT1_266
  (
    N744,
    N687
  );


  and
  AND2_267
  (
    N745,
    N228,
    N692
  );


  and
  AND2_268
  (
    N746,
    N237,
    N687
  );


  not
  NOT1_269
  (
    N747,
    N697
  );


  and
  AND2_270
  (
    N748,
    N228,
    N700
  );


  and
  AND2_271
  (
    N749,
    N237,
    N697
  );


  not
  NOT1_272
  (
    N750,
    N705
  );


  and
  AND2_273
  (
    N751,
    N228,
    N708
  );


  and
  AND2_274
  (
    N752,
    N237,
    N705
  );


  not
  NOT1_275
  (
    N753,
    N713
  );


  and
  AND2_276
  (
    N754,
    N228,
    N717
  );


  and
  AND2_277
  (
    N755,
    N237,
    N713
  );


  not
  NOT1_278
  (
    N756,
    N722
  );


  nor
  NOR2_279
  (
    N757,
    N727,
    N261
  );


  and
  AND2_280
  (
    N758,
    N727,
    N261
  );


  and
  AND2_281
  (
    N759,
    N228,
    N727
  );


  and
  AND2_282
  (
    N760,
    N237,
    N722
  );


  nand
  NAND2_283
  (
    N761,
    N644,
    N722
  );


  nand
  NAND2_284
  (
    N762,
    N635,
    N713
  );


  nand
  NAND3_285
  (
    N763,
    N635,
    N644,
    N722
  );


  nand
  NAND2_286
  (
    N764,
    N609,
    N687
  );


  nand
  NAND2_287
  (
    N765,
    N600,
    N678
  );


  nand
  NAND3_288
  (
    N766,
    N600,
    N609,
    N687
  );


  buf
  BUFF1_289
  (
    N767,
    N660
  );


  buf
  BUFF1_290
  (
    N768,
    N661
  );


  nor
  NOR2_291
  (
    N769,
    N736,
    N737
  );


  nor
  NOR2_292
  (
    N770,
    N739,
    N740
  );


  nor
  NOR2_293
  (
    N771,
    N742,
    N743
  );


  nor
  NOR2_294
  (
    N772,
    N745,
    N746
  );


  nand
  NAND4_295
  (
    N773,
    N750,
    N762,
    N763,
    N734
  );


  nor
  NOR2_296
  (
    N777,
    N748,
    N749
  );


  nand
  NAND3_297
  (
    N778,
    N753,
    N761,
    N733
  );


  nor
  NOR2_298
  (
    N781,
    N751,
    N752
  );


  nand
  NAND2_299
  (
    N782,
    N756,
    N732
  );


  nor
  NOR2_300
  (
    N785,
    N754,
    N755
  );


  nor
  NOR2_301
  (
    N786,
    N757,
    N758
  );


  nor
  NOR2_302
  (
    N787,
    N759,
    N760
  );


  nor
  NOR2_303
  (
    N788,
    N700,
    N773
  );


  and
  AND2_304
  (
    N789,
    N700,
    N773
  );


  nor
  NOR2_305
  (
    N790,
    N708,
    N778
  );


  and
  AND2_306
  (
    N791,
    N708,
    N778
  );


  nor
  NOR2_307
  (
    N792,
    N717,
    N782
  );


  and
  AND2_308
  (
    N793,
    N717,
    N782
  );


  and
  AND2_309
  (
    N794,
    N219,
    N786
  );


  nand
  NAND2_310
  (
    N795,
    N628,
    N773
  );


  nand
  NAND2_311
  (
    N796,
    N795,
    N747
  );


  nor
  NOR2_312
  (
    N802,
    N788,
    N789
  );


  nor
  NOR2_313
  (
    N803,
    N790,
    N791
  );


  nor
  NOR2_314
  (
    N804,
    N792,
    N793
  );


  nor
  NOR2_315
  (
    N805,
    N340,
    N794
  );


  nor
  NOR2_316
  (
    N806,
    N692,
    N796
  );


  and
  AND2_317
  (
    N807,
    N692,
    N796
  );


  and
  AND2_318
  (
    N808,
    N219,
    N802
  );


  and
  AND2_319
  (
    N809,
    N219,
    N803
  );


  and
  AND2_320
  (
    N810,
    N219,
    N804
  );


  nand
  NAND4_321
  (
    N811,
    N805,
    N787,
    N731,
    N529
  );


  nand
  NAND2_322
  (
    N812,
    N619,
    N796
  );


  nand
  NAND3_323
  (
    N813,
    N609,
    N619,
    N796
  );


  nand
  NAND4_324
  (
    N814,
    N600,
    N609,
    N619,
    N796
  );


  nand
  NAND4_325
  (
    N815,
    N738,
    N765,
    N766,
    N814
  );


  nand
  NAND3_326
  (
    N819,
    N741,
    N764,
    N813
  );


  nand
  NAND2_327
  (
    N822,
    N744,
    N812
  );


  nor
  NOR2_328
  (
    N825,
    N806,
    N807
  );


  nor
  NOR2_330
  (
    N827,
    N336,
    N809
  );


  not
  NOT1_332
  (
    N829,
    N811
  );


  nor
  NOR2_333
  (
    N830,
    N665,
    N815
  );


  and
  AND2_334
  (
    N831,
    N665,
    N815
  );


  nor
  NOR2_335
  (
    N832,
    N673,
    N819
  );


  and
  AND2_336
  (
    N833,
    N673,
    N819
  );


  nor
  NOR2_337
  (
    N834,
    N682,
    N822
  );


  and
  AND2_338
  (
    N835,
    N682,
    N822
  );


  and
  AND2_339
  (
    N836,
    N219,
    N825
  );


  nand
  NAND3_340
  (
    N837,
    N826,
    N777,
    N704
  );


  nand
  NAND4_341
  (
    N838,
    N827,
    N781,
    N712,
    N527
  );


  nand
  NAND4_342
  (
    N839,
    N828,
    N785,
    N721,
    N528
  );


  not
  NOT1_343
  (
    N840,
    N829
  );


  nand
  NAND2_344
  (
    N841,
    N815,
    N593
  );


  nor
  NOR2_345
  (
    N842,
    N830,
    N831
  );


  nor
  NOR2_346
  (
    N843,
    N832,
    N833
  );


  nor
  NOR2_347
  (
    N844,
    N834,
    N835
  );


  not
  NOT1_349
  (
    N846,
    N837
  );


  not
  NOT1_350
  (
    N847,
    N838
  );


  not
  NOT1_351
  (
    N848,
    N839
  );


  and
  AND2_352
  (
    N849,
    N735,
    N841
  );


  buf
  BUFF1_353
  (
    N850,
    N840
  );


  and
  AND2_354
  (
    N851,
    N219,
    N842
  );


  and
  AND2_355
  (
    N852,
    N219,
    N843
  );


  and
  AND2_356
  (
    N853,
    N219,
    N844
  );


  nand
  NAND3_357
  (
    N854,
    N845,
    N772,
    N696
  );


  not
  NOT1_358
  (
    N855,
    N846
  );


  not
  NOT1_360
  (
    N857,
    N848
  );


  not
  NOT1_361
  (
    N858,
    N849
  );


  nor
  NOR2_362
  (
    N859,
    N417,
    N851
  );


  nor
  NOR2_363
  (
    N860,
    N332,
    N852
  );


  nor
  NOR2_364
  (
    N861,
    N333,
    N853
  );


  not
  NOT1_365
  (
    N862,
    N854
  );


  buf
  BUFF1_366
  (
    N863,
    N855
  );


  buf
  BUFF1_367
  (
    N864,
    N856
  );


  buf
  BUFF1_368
  (
    N865,
    N857
  );


  buf
  BUFF1_369
  (
    N866,
    N858
  );


  nand
  NAND3_370
  (
    N867,
    N859,
    N769,
    N669
  );


  nand
  NAND3_371
  (
    N868,
    N860,
    N770,
    N677
  );


  nand
  NAND3_372
  (
    N869,
    N861,
    N771,
    N686
  );


  not
  NOT1_373
  (
    N870,
    N862
  );


  not
  NOT1_374
  (
    N871,
    N867
  );


  not
  NOT1_375
  (
    N872,
    N868
  );


  not
  NOT1_376
  (
    N873,
    N869
  );


  buf
  BUFF1_377
  (
    N874,
    N870
  );


  not
  NOT1_378
  (
    N875,
    N871
  );


  not
  NOT1_379
  (
    N876,
    N872
  );


  not
  NOT1_380
  (
    N877,
    N873
  );


  buf
  BUFF1_381
  (
    N878,
    N875
  );


  buf
  BUFF1_383
  (
    N880,
    N877
  );


  xor
  keyGate0
  (
    N644,
    keyWire0,
    keyInput0
  );


  or
  OR2_223
  (
    keyWire0,
    N577,
    N195
  );


  xor
  keyGate1
  (
    N517,
    keyWire1,
    keyInput1
  );


  and
  AND2_163
  (
    keyWire1,
    N126,
    N466
  );


  xnor
  keyGate2
  (
    N879,
    keyWire2,
    keyInput2
  );


  buf
  BUFF1_382
  (
    keyWire2,
    N876
  );


  xnor
  keyGate3
  (
    N524,
    keyWire3,
    keyInput3
  );


  and
  AND2_170
  (
    keyWire3,
    N451,
    N171
  );


  xor
  keyGate4
  (
    N826,
    keyWire4,
    keyInput4
  );


  nor
  NOR2_329
  (
    keyWire4,
    N335,
    N808
  );


  xor
  keyGate5
  (
    N845,
    keyWire5,
    keyInput5
  );


  nor
  NOR2_348
  (
    keyWire5,
    N334,
    N836
  );


  xor
  keyGate6
  (
    N423,
    keyWire6,
    keyInput6
  );


  buf
  BUFF1_109
  (
    keyWire6,
    N356
  );


  xor
  keyGate7
  (
    N659,
    keyWire7,
    keyInput7
  );


  and
  AND2_227
  (
    keyWire7,
    N246,
    N581
  );


  xor
  keyGate8
  (
    N539,
    keyWire8,
    keyInput8
  );


  nor
  NOR2_181
  (
    keyWire8,
    N318,
    N508
  );


  xnor
  keyGate9
  (
    N511,
    keyWire9,
    keyInput9
  );


  and
  AND2_157
  (
    keyWire9,
    N111,
    N466
  );


  xor
  keyGate10
  (
    N303,
    keyWire10,
    keyInput10
  );


  nand
  NAND2_22
  (
    keyWire10,
    N101,
    N106
  );


  xor
  keyGate11
  (
    N717,
    keyWire11,
    keyInput11
  );


  and
  AND2_249
  (
    keyWire11,
    N644,
    N641
  );


  xnor
  keyGate12
  (
    N590,
    keyWire12,
    keyInput12
  );


  nand
  NAND2_204
  (
    keyWire12,
    N553,
    N159
  );


  xor
  keyGate13
  (
    N279,
    keyWire13,
    keyInput13
  );


  nand
  NAND4_5
  (
    keyWire13,
    N1,
    N8,
    N51,
    N17
  );


  xor
  keyGate14
  (
    N355,
    keyWire14,
    keyInput14
  );


  nand
  NAND2_67
  (
    keyWire14,
    N89,
    N298
  );


  xnor
  keyGate15
  (
    N856,
    keyWire15,
    keyInput15
  );


  not
  NOT1_359
  (
    keyWire15,
    N847
  );


  xnor
  keyGate16
  (
    N389,
    keyWire16,
    keyInput16
  );


  buf
  BUFF1_80
  (
    keyWire16,
    N291
  );


  xor
  keyGate17
  (
    N305,
    keyWire17,
    keyInput17
  );


  nand
  NAND2_24
  (
    keyWire17,
    N111,
    N116
  );


  xnor
  keyGate18
  (
    N828,
    keyWire18,
    keyInput18
  );


  nor
  NOR2_331
  (
    keyWire18,
    N338,
    N810
  );


endmodule
